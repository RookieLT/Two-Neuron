`timescale 1ns/1ns
module tb_s1neuron;

//input 
reg [32*8-1 : 0] X;
reg [32*8-1 : 0] W;
//output
wire [31 : 0] H;
s1neuron #(8,32,12,20) dut (X,W,H);
initial begin
    X = 0;
    W = 0;
    #100;
    X = {32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000};
    W = {32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000};
end
endmodule