module row_weight #(parameter M=8,
                    parameter S=8,
                    parameter n=32,
                    parameter addrwidth=2)(
        input [addrwidth:0] addr,
        output [M*n-1 : 0] W
);

    reg [M*n-1 : 0] weight[S:0] ;
    initial begin
        
        weight[0]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[1]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[2]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[3]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[4]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[5]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[6]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[7]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[8]='b0;
    end

assign W = weight[addr];

endmodule