`timescale 1ns/1ns
module tb_s2neuron;
//input 
reg [31 : 0] H;
reg [32*8-1 : 0] W;
reg finished;
//output
wire [255 : 0] Y;
s2neuron #(8,8,32,12,20) dut (H,W,finished,Y);
initial begin
    H = 32'b0000_0000_0001_0000_0000_0000_0000_0000;
    W = {32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000};
    #20;
    H = 32'b0000_0000_0000_1000_0000_0000_0000_0000;
    W = {32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000};
    finished =1;
end
endmodule