module row_weight #(parameter M=8,
                    parameter S=8,
                    parameter n=32)(
        input [2:0] addr,
        output [M*n-1 : 0] W
);

    reg [M*n-1 : 0] weight[S-1:0] ;
    initial begin
        weight[0]={32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[1]={32'h00001000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[2]={32'h00010100,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[3]={32'h00010010,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[4]={32'h00010001,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[5]={32'h00010010,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[6]={32'h00010100,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[7]={32'h00011000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
    end

assign W = weight[addr];

endmodule