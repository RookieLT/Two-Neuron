`timescale 1ns/1ns
module tb_rmac;

//input
reg [31:0] W,X;
reg finished;
//output
wire [31:0] sum;

initial begin
    finished=0;
    W=32'b0000_0000_0001_0000_0000_0000_0000_0000;
    X=32'b0000_0000_0001_0000_0000_0000_0000_0000;
    #10;
    W=32'b0000_0000_0000_1000_0000_0000_0000_0000;
    X=32'b0000_0000_0001_0000_0000_0000_0000_0000;
    #10;
    W=32'b0000_0000_0000_1100_0000_0000_0000_0000;
    X=32'b0000_0000_0001_0000_0000_0000_0000_0000;
    finished = 1;
end

rmac #(8,32,12,20) dut(W,X,finished,sum); 
endmodule