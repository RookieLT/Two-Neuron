module column_weight #(parameter N=8,
                    parameter S=8,
                    parameter n=32,
                    parameter addrwidth=2)(
        input [addrwidth:0] addr,
        output [N*n-1 : 0] W
);


    reg [N*n-1 : 0] weight[S:0] ;
    initial begin
        /*weight[0]={32'h00011000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[1]={32'h00010100,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[2]={32'h00010010,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[3]={32'h00010001,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[4]={32'h00010010,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[5]={32'h00010100,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[6]={32'h00011000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};
        weight[7]={32'h00010100,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000,32'h00010000};*/
        /*weight[0]={16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066};
        weight[1]={16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066};
        weight[2]={16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066,16'h0066};
        weight[3]={16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066};
        weight[4]={16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066};
        weight[5]={16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066,16'h8066};
        weight[6]={16'h0200,16'h0200,16'h0200,16'h0200,16'h0200,16'h0200,16'h0200,16'h0200};
        weight[7]={16'h0200,16'h0200,16'h0200,16'h0200,16'h0200,16'h0200,16'h0200,16'h0200};*/
        weight[0]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[1]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        weight[2]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[3]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        weight[4]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[5]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        weight[6]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[7]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        weight[8]='b0;
    end

assign W = weight[addr];
endmodule