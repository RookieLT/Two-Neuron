`timescale 1ns/1ns
module tb_top;

//input
reg clk,reset;
reg [255:0] X;
//output
wire [255:0] Y;
top #(8,8,8,32,12,20) TP(clk,reset,X,Y);
initial begin
    clk=0;
    forever begin
        #10 clk=!clk;
    end
end
initial begin
    reset =1;
    #20;
    reset=0;
    #300;
    reset =1;
    #20;
    reset=0;
end
initial begin
    X =  {32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000,
        32'b0000_0000_0001_0000_0000_0000_0000_0000};
end
endmodule