module mlp_ctrl#(parameter M=784,
                parameter N=512,
                parameter S=512,
                parameter K=16)(
                input clk,rst,
                input 
                );